module tb_simon32x64()
endmodule

